
`timescale 1ns / 1ps

module fifo_top #(
    parameter DATASIZE = 8,             // Data width. This is the size of our data to be read of written which is of 8-bits
    parameter ADDRSIZE = 4              // Address width. 2^4 = 16. Hence the depth of our FIFO is 16. This address will be used to map to the pointer 0 - 15
)(
    output logic [DATASIZE-1:0] rdata,  // data that would be read out from FIFO
    output logic wfull,  // FIFO is full indication so cannot write anymore
    output logic rempty, // FIFO is empty so nothing to read 
    output logic walmost_full, // Write side 3/4th full
    output logic ralmost_empty, // read side 3/4th full
    input logic [DATASIZE-1:0] wdata, // data that should be written into FIFO
    input logic winc, wclk, wrst_n, //winc is our write enable, wclk the clk for write doman and wrst_n is our active low reset for write domain
    input logic rinc, rclk, rrst_n //rinc is the read enable, rclk is the clk for read domain and rrst_n is our active low reset for read domain
);

    logic [ADDRSIZE-1:0] waddr;  // The write address used to index memory on wclk
    logic [ADDRSIZE-1:0] raddr; // The read address used to index memory on rclk
    logic [ADDRSIZE:0] wptr; // The write pointer in gray code generated by the write side. This will be sent across the clock domain into the read domain
    logic [ADDRSIZE:0] rptr; // The read pointer in gray code generated by the read side. This will be sent across the clock domain into the write domain
    logic [ADDRSIZE:0] wq2_rptr; // This is the read pointer after the 2-FF synchronization into the write clock domain
    logic [ADDRSIZE:0] rq2_wptr; // This is the write pointer after the 2-FF synchronization into the read clock domain

    fifo_sync_r2w sync_r2w (            // Instantiation of synchronizer from read to write domain
        .*                              // This module brings the read pointer rptr into the write clock domain
    );                                  // .* connects all signals with the same name

    fifo_sync_w2r sync_w2r (            // Instantiation of synchronizer from write to read domain
        .*                              // This module brings the write pointer wptr into the read clock domain
    );                                  // .* connects all signals with the same name 

    fifo_memory #(                      // Our FIFO memory module
        .DATASIZE(DATASIZE),            // 8-bit data size
        .ADDRSIZE(ADDRSIZE)             // 4-bit address representation
    ) fifomem (
        .rdata(rdata),                  // All signals connected respectively to the top
        .wdata(wdata),
        .waddr(waddr),
        .raddr(raddr),
        .wclken(winc),
        .wfull(wfull),
        .wclk(wclk)
    );

    fifo_read #(ADDRSIZE) rptr_empty (  // Read side controller module
        .*
    );

    fifo_write #(ADDRSIZE) wptr_full (  // Write side controller module
        .*
    );

endmodule

